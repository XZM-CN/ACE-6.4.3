128 path=ACE_wrappers/performance-tests/Server_Concurrency/Queue_Based_Workers/GNUmakefile.Svr_Conc_Queue_Based_Workers_RTCorba
30 mtime=1492674765.548638377
30 atime=1492675753.319045631
30 ctime=1492675751.411048611
